module fetch_tb;


initial
begin
  $display("CPU | Fetch		testbench");

  $finish;
end

endmodule
